module mem_arb
